module srff_tb;
  reg clk, S, R;
  wire Q;

  srff dut(.clk(clk), .S(S), .R(R), .Q(Q));

  initial begin
    clk = 0;
    forever #10 clk = ~clk;
  end

  initial begin
    S = 0; R = 0;
    #100 S = 1; R = 0;
    #100 S = 0; R = 0;
    #100 S = 0; R = 1;
    #100 S = 1; R = 1;
    #100 S = 0; R = 0;
  end
endmodule
